* /Users/peterkinget/Library/Mobile Documents/com~apple~CloudDocs/Work/MOBIUS/GitHub/adding_connections_to_bitstream/MobiusCADFlow/LTspice/examples/library 3stage_RO tsmc025_public/7stage_RO_schematic.asc
XX4 BUS05 BUS06 BUS09 dp_nmos_1x_a
XX5 BUS05 BUS06 BUS09 dp_nmos_1x_b
XX2 BUS06 BUS07 cs_nmos_4x_a
XX6 BUS03 BUS04 BUS09 BUS09 dp_nmos_4x_a
XX7 BUS04 BUS05 BUS09 BUS09 dp_nmos_4x_b
XX9 BUS07 BUS06 cs_pmos_4x_a
XX10 BUS01 BUS07 cs_pmos_4x_b
XX3 BUS07 BUS01 cs_nmos_4x_b
XX13 BUS04 BUS03 BUS10 BUS10 dp_pmos_4x_a
XX14 BUS05 BUS04 BUS10 BUS10 dp_pmos_4x_b
XX15 BUS06 BUS05 BUS10 dp_pmos_1x_b
XX16 BUS06 BUS05 BUS10 dp_pmos_1x_a
XX17 BUS02 BUS02 BUS03 inverter_a
XX18 BUS01 BUS01 BUS02 inverter_b
XX21 BUS10 chip_vdd
XX22 BUS09 chip_vss
V2 VDD 0 {VDD}
I1 BUS07 BUS09 PWL(0 0 10n 1m 20n 0)
C1 BUS02 BUS09 {Cpar}
C2 BUS03 BUS09 {Cpar}
C3 BUS04 BUS09 {Cpar}
C4 BUS05 BUS09 {Cpar}
C5 BUS06 BUS09 {Cpar}
C6 BUS07 BUS09 {Cpar}
C7 BUS01 BUS09 {Cpar}

* block symbol definitions
.subckt dp_nmos_1x_a gate drain source
XM1 drain gate source 0 NMOS_mobius m=1
.ends dp_nmos_1x_a

.subckt dp_nmos_1x_b gate drain source
XM1 drain gate source 0 NMOS_mobius m=1
.ends dp_nmos_1x_b

.subckt cs_nmos_4x_a gate drain
XM1 drain gate 0 0 NMOS_mobius m=4
.ends cs_nmos_4x_a

.subckt dp_nmos_4x_a gate drain source substrate
XM1 drain gate source substrate NMOS_mobius m=4
.ends dp_nmos_4x_a

.subckt dp_nmos_4x_b gate drain source substrate
XM1 drain gate source substrate NMOS_mobius m=4
.ends dp_nmos_4x_b

.subckt cs_pmos_4x_a drain gate
XM1 drain gate VDD VDD PMOS_mobius m=4
.ends cs_pmos_4x_a

.subckt cs_pmos_4x_b drain gate
XM1 drain gate VDD VDD PMOS_mobius m=4
.ends cs_pmos_4x_b

.subckt cs_nmos_4x_b gate drain
XM1 drain gate 0 0 NMOS_mobius m=4
.ends cs_nmos_4x_b

.subckt dp_pmos_4x_a drain gate source nwell
XM1 drain gate source nwell PMOS_mobius m=4
.ends dp_pmos_4x_a

.subckt dp_pmos_4x_b drain gate source nwell
XM1 drain gate source nwell PMOS_mobius m=4
.ends dp_pmos_4x_b

.subckt dp_pmos_1x_b drain gate source
XM1 drain gate source VDD PMOS_mobius m=1
.ends dp_pmos_1x_b

.subckt dp_pmos_1x_a drain gate source
XM1 drain gate source VDD PMOS_mobius m=1
.ends dp_pmos_1x_a

.subckt inverter_a inn inp out
XM1 out inn 0 0 NMOS_mobius m=16
XM2 out inp VDD VDD PMOS_mobius m=16
.ends inverter_a

.subckt inverter_b inn inp out
XM1 out inn 0 0 NMOS_mobius m=16
XM2 out inp VDD VDD PMOS_mobius m=16
.ends inverter_b

.subckt chip_vdd chip_vdd
R1 chip_vdd VDD .000001
.ends chip_vdd

.subckt chip_vss chip_vss
R1 chip_vss 0 0.000001
.ends chip_vss

* Note: Do not connect a BUS directly to VDD or VSS even with a jumper. \nUse the Chip_VDD and Chip_VSS.
* Seven Stage Ring Oscillator 16-16-4-4-2-4-4\n7stage_RO
.global VDD
.param VDD = 2.5
.inc transistor_models_tsmc025_public.inc
.tran 10u
.meas tran zc1 find time when v(bus01) = 1.25 rise=20
.meas tran zc2 find time when v(bus01) = 1.25 rise=21
.meas tran freq param 1/(zc2-zc1)
.param Cpar=200p
* Models and Global Parameters
* Measurements
* Circuit Parameters
* Simulation Command
* Note: Do not connect a BUS directly to VDD or VSS even with a jumper. Use the Chip_VDD and Chip_VSS.
.backanno
.end
