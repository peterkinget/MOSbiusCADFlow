* /Users/peterkinget/Library/Mobile Documents/com~apple~CloudDocs/Work/MOBIUS/LTSpice_working_area/library Miller OTA pMOS tsmc025_public/Miller_OTA_pin.asc
XX1 BUS02 BUS03 nmos_currentmirror
XX2 BUS03 BUS04 cs_nmos_4x_a
XX6 BUS03 BUS04 BUS09 BUS09 dp_nmos_4x_a
XX7 BUS03 BUS04 BUS09 BUS09 dp_nmos_4x_b
V1 VDD 0 {VDD}
XX12 N001 NC_01 BUS01 NC_02 NC_03 BUS04 pmos_currentmirror_array
XX3 BUS03 BUS04 cs_nmos_4x_b
XX13 BUS02 N002 BUS01 BUS01 dp_pmos_4x_a
XX14 BUS03 vinp BUS01 BUS01 dp_pmos_4x_b
XX22 BUS09 chip_vss
I1 N001 0 {IBIAS}
V2 vinp 0 {VDD/2} AC 1
C1 BUS04 0 {Cload}
C2 N002 0 {Clarge}
L1 N002 N004 {Llarge}
E1 N004 0 BUS04 0 1
C3 BUS04 N003 {Ccomp}
R1 N003 BUS03 {Rcomp}

* block symbol definitions
.subckt nmos_currentmirror in out
XM1 in in 0 0 NMOS_mobius m=1
XM2 out in 0 0 NMOS_mobius m=1
.ends nmos_currentmirror

.subckt cs_nmos_4x_a gate drain
XM1 drain gate 0 0 NMOS_mobius m=4
.ends cs_nmos_4x_a

.subckt dp_nmos_4x_a gate drain source substrate
XM1 drain gate source substrate NMOS_mobius m=4
.ends dp_nmos_4x_a

.subckt dp_nmos_4x_b gate drain source substrate
XM1 drain gate source substrate NMOS_mobius m=4
.ends dp_nmos_4x_b

.subckt pmos_currentmirror_array in out1 out2 out4 out8 out16
XM1 in in VDD VDD PMOS_mobius m=1
XM2 out1 in VDD VDD PMOS_mobius m=1
XM3 out2 in VDD VDD PMOS_mobius m=2
XM4 out4 in VDD VDD PMOS_mobius m=4
XM5 out8 in VDD VDD PMOS_mobius m=8
XM6 out16 in VDD VDD PMOS_mobius m=16
.ends pmos_currentmirror_array

.subckt cs_nmos_4x_b gate drain
XM1 drain gate 0 0 NMOS_mobius m=4
.ends cs_nmos_4x_b

.subckt dp_pmos_4x_a drain gate source nwell
XM1 drain gate source nwell PMOS_mobius m=4
.ends dp_pmos_4x_a

.subckt dp_pmos_4x_b drain gate source nwell
XM1 drain gate source nwell PMOS_mobius m=4
.ends dp_pmos_4x_b

.subckt chip_vss chip_vss
R1 chip_vss 0 0.000001
.ends chip_vss

.global VDD
.param VDD = 2.5
.inc transistor_models_tsmc025_public.inc
*.step param Ccomp list 100f 100p 200p 400p
*.step param Rcomp list 0.001 200
*.ac dec 50 1 1e9
.op
* Note: Do not connect a BUS directly to VDD or VSS even with a jumper. \nUse the Chip_VDD and Chip_VSS.
.param IBIAS = 100u Cload = 200p Ccomp=120p Rcomp=200
.param Clarge = 10 Llarge = 10
.backanno
.end
