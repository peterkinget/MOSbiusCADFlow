* /Users/peterkinget/Library/Mobile Documents/com~apple~CloudDocs/Work/MOBIUS/GitHub/adding_connections_to_bitstream/MobiusCADFlow/LTspice/examples/library 3stage_RO tsmc025_public/3stage_RO_8x_schematic.asc
XX6 BUS03 BUS01 BUS10 BUS10 dp_nmos_4x_a
XX7 BUS03 BUS01 BUS10 BUS10 dp_nmos_4x_b
V1 VDD 0 {VDD}
XX13 BUS01 BUS03 BUS09 BUS09 dp_pmos_4x_a
XX14 BUS01 BUS03 BUS09 BUS09 dp_pmos_4x_b
XX17 BUS02 BUS02 BUS03 inverter_a
XX18 BUS01 BUS01 BUS02 inverter_b
I1 BUS01 BUS10 PWL(0 0 10n 1m 20n 0)
C1 BUS02 BUS10 {Cpar}
C2 BUS03 BUS10 {Cpar}
C3 BUS01 BUS10 {Cpar}
XX1 BUS09 chip_vdd
XX2 BUS10 chip_vss

* block symbol definitions
.subckt dp_nmos_4x_a gate drain source substrate
XM1 drain gate source substrate NMOS_mobius m=4
.ends dp_nmos_4x_a

.subckt dp_nmos_4x_b gate drain source substrate
XM1 drain gate source substrate NMOS_mobius m=4
.ends dp_nmos_4x_b

.subckt dp_pmos_4x_a drain gate source nwell
XM1 drain gate source nwell PMOS_mobius m=4
.ends dp_pmos_4x_a

.subckt dp_pmos_4x_b drain gate source nwell
XM1 drain gate source nwell PMOS_mobius m=4
.ends dp_pmos_4x_b

.subckt inverter_a inn inp out
XM1 out inn 0 0 NMOS_mobius m=16
XM2 out inp VDD VDD PMOS_mobius m=16
.ends inverter_a

.subckt inverter_b inn inp out
XM1 out inn 0 0 NMOS_mobius m=16
XM2 out inp VDD VDD PMOS_mobius m=16
.ends inverter_b

.subckt chip_vdd chip_vdd
R1 chip_vdd VDD .000001
.ends chip_vdd

.subckt chip_vss chip_vss
R1 chip_vss 0 0.000001
.ends chip_vss

.global VDD
.param VDD = 2.5
.inc transistor_models_tsmc025_public.inc
.tran 5u
.meas tran zc1 find time when v(bus01) = 1.25 rise=20
.meas tran zc2 find time when v(bus01) = 1.25 rise=21
.meas tran freq param 1/(zc2-zc1)
.param Cpar=200p
* Models and Global Parameters
* Measurements
* Circuit Parameters
* Simulation Command
* Three Stage Ring Oscillator 16-16-8\n3stage_RO_8x
* for startup
* Note: Do not connect a BUS directly to VDD or VSS even with a jumper. Use the Chip_VDD and Chip_VSS.
.backanno
.end
